module rv_go_iiiii (
	ports
);
	
endmodule